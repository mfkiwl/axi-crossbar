// distributed under the mit license
// https://opensource.org/licenses/mit-license.php

///////////////////////////////////////////////////////////////////////////////
//
// AXI4 crossbar top level, instanciating the global infrastructure of the
// core. All the master and slave interfaces are instanciated here.
//
///////////////////////////////////////////////////////////////////////////////

`timescale 1 ns / 1 ps
`default_nettype none

module axi_crossbar_top

    #(
        // Address bus width
        parameter ADDR_W = 8,
        // AXI ID width
        parameter AXI_ID_W = 8,
        // AXI4 data width
        parameter AXI_DATA_W = 8
    )(
        // Interconnect global interface
        input  logic                      aclk,
        input  logic                      aresetn,
        input  logic                      srst,
        // Master 0 interface
        input  logic                      mst0_awvalid,
        output logic                      mst0_awready,
        input  logic [ADDR_W        -1:0] mst0_awaddr,
        input  logic [8             -1:0] mst0_awlen,
        input  logic [3             -1:0] mst0_awsize,
        input  logic [2             -1:0] mst0_awburst,
        input  logic [2             -1:0] mst0_awlock,
        input  logic [4             -1:0] mst0_awcache,
        input  logic [3             -1:0] mst0_awprot,
        input  logic [4             -1:0] mst0_awqos,
        input  logic [4             -1:0] mst0_awregion,
        input  logic [AXI_ID_W      -1:0] mst0_awid,
        input  logic                      mst0_wvalid,
        output logic                      mst0_wready,
        input  logic                      mst0_wlast,
        input  logic [AXI_DATA_W    -1:0] mst0_wdata,
        input  logic [AXI_DATA_W/8  -1:0] mst0_wstrb,
        output logic                      mst0_bvalid,
        input  logic                      mst0_bready,
        output logic [AXI_ID_W      -1:0] mst0_bid,
        output logic [2             -1:0] mst0_bresp,
        input  logic                      mst0_arvalid,
        output logic                      mst0_arready,
        input  logic [ADDR_W        -1:0] mst0_araddr,
        input  logic [8             -1:0] mst0_arlen,
        input  logic [3             -1:0] mst0_arsize,
        input  logic [2             -1:0] mst0_arburst,
        input  logic [2             -1:0] mst0_arlock,
        input  logic [4             -1:0] mst0_arcache,
        input  logic [3             -1:0] mst0_arprot,
        input  logic [4             -1:0] mst0_arqos,
        input  logic [4             -1:0] mst0_arregion,
        input  logic [AXI_ID_W      -1:0] mst0_arid,
        output logic                      mst0_rvalid,
        input  logic                      mst0_rready,
        output logic [AXI_ID_W      -1:0] mst0_rid,
        output logic [2             -1:0] mst0_rresp,
        output logic [AXI_DATA_W    -1:0] mst0_rdata,
        output logic                      mst0_rlast,
        // Master 1 interface
        input  logic                      mst1_awvalid,
        output logic                      mst1_awready,
        input  logic [ADDR_W        -1:0] mst1_awaddr,
        input  logic [8             -1:0] mst1_awlen,
        input  logic [3             -1:0] mst1_awsize,
        input  logic [2             -1:0] mst1_awburst,
        input  logic [2             -1:0] mst1_awlock,
        input  logic [4             -1:0] mst1_awcache,
        input  logic [3             -1:0] mst1_awprot,
        input  logic [4             -1:0] mst1_awqos,
        input  logic [4             -1:0] mst1_awregion,
        input  logic [AXI_ID_W      -1:0] mst1_awid,
        input  logic                      mst1_wvalid,
        output logic                      mst1_wready,
        input  logic                      mst1_wlast,
        input  logic [AXI_DATA_W    -1:0] mst1_wdata,
        input  logic [AXI_DATA_W/8  -1:0] mst1_wstrb,
        output logic                      mst1_bvalid,
        input  logic                      mst1_bready,
        output logic [AXI_ID_W      -1:0] mst1_bid,
        output logic [2             -1:0] mst1_bresp,
        input  logic                      mst1_arvalid,
        output logic                      mst1_arready,
        input  logic [ADDR_W        -1:0] mst1_araddr,
        input  logic [8             -1:0] mst1_arlen,
        input  logic [3             -1:0] mst1_arsize,
        input  logic [2             -1:0] mst1_arburst,
        input  logic [2             -1:0] mst1_arlock,
        input  logic [4             -1:0] mst1_arcache,
        input  logic [3             -1:0] mst1_arprot,
        input  logic [4             -1:0] mst1_arqos,
        input  logic [4             -1:0] mst1_arregion,
        input  logic [AXI_ID_W      -1:0] mst1_arid,
        output logic                      mst1_rvalid,
        input  logic                      mst1_rready,
        output logic [AXI_ID_W      -1:0] mst1_rid,
        output logic [2             -1:0] mst1_rresp,
        output logic [AXI_DATA_W    -1:0] mst1_rdata,
        output logic                      mst1_rlast,
        // Master 1 interface
        input  logic                      mst2_awvalid,
        output logic                      mst2_awready,
        input  logic [ADDR_W        -1:0] mst2_awaddr,
        input  logic [8             -1:0] mst2_awlen,
        input  logic [3             -1:0] mst2_awsize,
        input  logic [2             -1:0] mst2_awburst,
        input  logic [2             -1:0] mst2_awlock,
        input  logic [4             -1:0] mst2_awcache,
        input  logic [3             -1:0] mst2_awprot,
        input  logic [4             -1:0] mst2_awqos,
        input  logic [4             -1:0] mst2_awregion,
        input  logic [AXI_ID_W      -1:0] mst2_awid,
        input  logic                      mst2_wvalid,
        output logic                      mst2_wready,
        input  logic                      mst2_wlast,
        input  logic [AXI_DATA_W    -1:0] mst2_wdata,
        input  logic [AXI_DATA_W/8  -1:0] mst2_wstrb,
        output logic                      mst2_bvalid,
        input  logic                      mst2_bready,
        output logic [AXI_ID_W      -1:0] mst2_bid,
        output logic [2             -1:0] mst2_bresp,
        input  logic                      mst2_arvalid,
        output logic                      mst2_arready,
        input  logic [ADDR_W        -1:0] mst2_araddr,
        input  logic [8             -1:0] mst2_arlen,
        input  logic [3             -1:0] mst2_arsize,
        input  logic [2             -1:0] mst2_arburst,
        input  logic [2             -1:0] mst2_arlock,
        input  logic [4             -1:0] mst2_arcache,
        input  logic [3             -1:0] mst2_arprot,
        input  logic [4             -1:0] mst2_arqos,
        input  logic [4             -1:0] mst2_arregion,
        input  logic [AXI_ID_W      -1:0] mst2_arid,
        output logic                      mst2_rvalid,
        input  logic                      mst2_rready,
        output logic [AXI_ID_W      -1:0] mst2_rid,
        output logic [2             -1:0] mst2_rresp,
        output logic [AXI_DATA_W    -1:0] mst2_rdata,
        output logic                      mst2_rlast,
        // Master 1 interface
        input  logic                      mst3_awvalid,
        output logic                      mst3_awready,
        input  logic [ADDR_W        -1:0] mst3_awaddr,
        input  logic [8             -1:0] mst3_awlen,
        input  logic [3             -1:0] mst3_awsize,
        input  logic [2             -1:0] mst3_awburst,
        input  logic [2             -1:0] mst3_awlock,
        input  logic [4             -1:0] mst3_awcache,
        input  logic [3             -1:0] mst3_awprot,
        input  logic [4             -1:0] mst3_awqos,
        input  logic [4             -1:0] mst3_awregion,
        input  logic [AXI_ID_W      -1:0] mst3_awid,
        input  logic                      mst3_wvalid,
        output logic                      mst3_wready,
        input  logic                      mst3_wlast,
        input  logic [AXI_DATA_W    -1:0] mst3_wdata,
        input  logic [AXI_DATA_W/8  -1:0] mst3_wstrb,
        output logic                      mst3_bvalid,
        input  logic                      mst3_bready,
        output logic [AXI_ID_W      -1:0] mst3_bid,
        output logic [2             -1:0] mst3_bresp,
        input  logic                      mst3_arvalid,
        output logic                      mst3_arready,
        input  logic [ADDR_W        -1:0] mst3_araddr,
        input  logic [8             -1:0] mst3_arlen,
        input  logic [3             -1:0] mst3_arsize,
        input  logic [2             -1:0] mst3_arburst,
        input  logic [2             -1:0] mst3_arlock,
        input  logic [4             -1:0] mst3_arcache,
        input  logic [3             -1:0] mst3_arprot,
        input  logic [4             -1:0] mst3_arqos,
        input  logic [4             -1:0] mst3_arregion,
        input  logic [AXI_ID_W      -1:0] mst3_arid,
        output logic                      mst3_rvalid,
        input  logic                      mst3_rready,
        output logic [AXI_ID_W      -1:0] mst3_rid,
        output logic [2             -1:0] mst3_rresp,
        output logic [AXI_DATA_W    -1:0] mst3_rdata,
        output logic                      mst3_rlast,
        // Slave 0 interface
        output logic                      slv0_awvalid,
        input  logic                      slv0_awready,
        output logic [ADDR_W        -1:0] slv0_awaddr,
        output logic [8             -1:0] slv0_awlen,
        output logic [3             -1:0] slv0_awsize,
        output logic [2             -1:0] slv0_awburst,
        output logic [2             -1:0] slv0_awlock,
        output logic [4             -1:0] slv0_awcache,
        output logic [3             -1:0] slv0_awprot,
        output logic [4             -1:0] slv0_awqos,
        output logic [4             -1:0] slv0_awregion,
        output logic [AXI_ID_W      -1:0] slv0_awid,
        output logic                      slv0_wvalid,
        input  logic                      slv0_wready,
        input  logic                      slv0_wlast,
        output logic [AXI_DATA_W    -1:0] slv0_wdata,
        output logic [AXI_DATA_W/8  -1:0] slv0_wstrb,
        input  logic                      slv0_bvalid,
        output logic                      slv0_bready,
        input  logic [AXI_ID_W      -1:0] slv0_bid,
        input  logic [2             -1:0] slv0_bresp,
        output logic                      slv0_arvalid,
        input  logic                      slv0_arready,
        output logic [ADDR_W        -1:0] slv0_araddr,
        output logic [8             -1:0] slv0_arlen,
        output logic [3             -1:0] slv0_arsize,
        output logic [2             -1:0] slv0_arburst,
        output logic [2             -1:0] slv0_arlock,
        output logic [4             -1:0] slv0_arcache,
        output logic [3             -1:0] slv0_arprot,
        output logic [4             -1:0] slv0_arqos,
        output logic [4             -1:0] slv0_arregion,
        output logic [AXI_ID_W      -1:0] slv0_arid,
        input  logic                      slv0_rvalid,
        output logic                      slv0_rready,
        input  logic [AXI_ID_W      -1:0] slv0_rid,
        input  logic [2             -1:0] slv0_rresp,
        input  logic [AXI_DATA_W    -1:0] slv0_rdata,
        input  logic                      slv0_rlast,
        // Slave 1 interface
        output logic                      slv1_awvalid,
        input  logic                      slv1_awready,
        output logic [ADDR_W        -1:0] slv1_awaddr,
        output logic [8             -1:0] slv1_awlen,
        output logic [3             -1:0] slv1_awsize,
        output logic [2             -1:0] slv1_awburst,
        output logic [2             -1:0] slv1_awlock,
        output logic [4             -1:0] slv1_awcache,
        output logic [3             -1:0] slv1_awprot,
        output logic [4             -1:0] slv1_awqos,
        output logic [4             -1:0] slv1_awregion,
        output logic [AXI_ID_W      -1:0] slv1_awid,
        output logic                      slv1_wvalid,
        input  logic                      slv1_wready,
        input  logic                      slv1_wlast,
        output logic [AXI_DATA_W    -1:0] slv1_wdata,
        output logic [AXI_DATA_W/8  -1:0] slv1_wstrb,
        input  logic                      slv1_bvalid,
        output logic                      slv1_bready,
        input  logic [AXI_ID_W      -1:0] slv1_bid,
        input  logic [2             -1:0] slv1_bresp,
        output logic                      slv1_arvalid,
        input  logic                      slv1_arready,
        output logic [ADDR_W        -1:0] slv1_araddr,
        output logic [8             -1:0] slv1_arlen,
        output logic [3             -1:0] slv1_arsize,
        output logic [2             -1:0] slv1_arburst,
        output logic [2             -1:0] slv1_arlock,
        output logic [4             -1:0] slv1_arcache,
        output logic [3             -1:0] slv1_arprot,
        output logic [4             -1:0] slv1_arqos,
        output logic [4             -1:0] slv1_arregion,
        output logic [AXI_ID_W      -1:0] slv1_arid,
        input  logic                      slv1_rvalid,
        output logic                      slv1_rready,
        input  logic [AXI_ID_W      -1:0] slv1_rid,
        input  logic [2             -1:0] slv1_rresp,
        input  logic [AXI_DATA_W    -1:0] slv1_rdata,
        input  logic                      slv1_rlast,
        // Slave 2 interface
        output logic                      slv2_awvalid,
        input  logic                      slv2_awready,
        output logic [ADDR_W        -1:0] slv2_awaddr,
        output logic [8             -1:0] slv2_awlen,
        output logic [3             -1:0] slv2_awsize,
        output logic [2             -1:0] slv2_awburst,
        output logic [2             -1:0] slv2_awlock,
        output logic [4             -1:0] slv2_awcache,
        output logic [3             -1:0] slv2_awprot,
        output logic [4             -1:0] slv2_awqos,
        output logic [4             -1:0] slv2_awregion,
        output logic [AXI_ID_W      -1:0] slv2_awid,
        output logic                      slv2_wvalid,
        input  logic                      slv2_wready,
        input  logic                      slv2_wlast,
        output logic [AXI_DATA_W    -1:0] slv2_wdata,
        output logic [AXI_DATA_W/8  -1:0] slv2_wstrb,
        input  logic                      slv2_bvalid,
        output logic                      slv2_bready,
        input  logic [AXI_ID_W      -1:0] slv2_bid,
        input  logic [2             -1:0] slv2_bresp,
        output logic                      slv2_arvalid,
        input  logic                      slv2_arready,
        output logic [ADDR_W        -1:0] slv2_araddr,
        output logic [8             -1:0] slv2_arlen,
        output logic [3             -1:0] slv2_arsize,
        output logic [2             -1:0] slv2_arburst,
        output logic [2             -1:0] slv2_arlock,
        output logic [4             -1:0] slv2_arcache,
        output logic [3             -1:0] slv2_arprot,
        output logic [4             -1:0] slv2_arqos,
        output logic [4             -1:0] slv2_arregion,
        output logic [AXI_ID_W      -1:0] slv2_arid,
        input  logic                      slv2_rvalid,
        output logic                      slv2_rready,
        input  logic [AXI_ID_W      -1:0] slv2_rid,
        input  logic [2             -1:0] slv2_rresp,
        input  logic [AXI_DATA_W    -1:0] slv2_rdata,
        input  logic                      slv2_rlast,
        // Slave 3 interface
        output logic                      slv3_awvalid,
        input  logic                      slv3_awready,
        output logic [ADDR_W        -1:0] slv3_awaddr,
        output logic [8             -1:0] slv3_awlen,
        output logic [3             -1:0] slv3_awsize,
        output logic [2             -1:0] slv3_awburst,
        output logic [2             -1:0] slv3_awlock,
        output logic [4             -1:0] slv3_awcache,
        output logic [3             -1:0] slv3_awprot,
        output logic [4             -1:0] slv3_awqos,
        output logic [4             -1:0] slv3_awregion,
        output logic [AXI_ID_W      -1:0] slv3_awid,
        output logic                      slv3_wvalid,
        input  logic                      slv3_wready,
        input  logic                      slv3_wlast,
        output logic [AXI_DATA_W    -1:0] slv3_wdata,
        output logic [AXI_DATA_W/8  -1:0] slv3_wstrb,
        input  logic                      slv3_bvalid,
        output logic                      slv3_bready,
        input  logic [AXI_ID_W      -1:0] slv3_bid,
        input  logic [2             -1:0] slv3_bresp,
        output logic                      slv3_arvalid,
        input  logic                      slv3_arready,
        output logic [ADDR_W        -1:0] slv3_araddr,
        output logic [8             -1:0] slv3_arlen,
        output logic [3             -1:0] slv3_arsize,
        output logic [2             -1:0] slv3_arburst,
        output logic [2             -1:0] slv3_arlock,
        output logic [4             -1:0] slv3_arcache,
        output logic [3             -1:0] slv3_arprot,
        output logic [4             -1:0] slv3_arqos,
        output logic [4             -1:0] slv3_arregion,
        output logic [AXI_ID_W      -1:0] slv3_arid,
        input  logic                      slv3_rvalid,
        output logic                      slv3_rready,
        input  logic [AXI_ID_W      -1:0] slv3_rid,
        input  logic [2             -1:0] slv3_rresp,
        input  logic [AXI_DATA_W    -1:0] slv3_rdata,
        input  logic                      slv3_rlast
    );


endmodule

`resetall

